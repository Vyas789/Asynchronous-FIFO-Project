`define DATA 8
`define no_of_trans 20
`define ADDR 4
`define WIDTH 8
      
