//`include "uvm_macros.svh"
package async_fifo_pkg;
    
    `include "uvm_macros.svh"
	import uvm_pkg::*;
    `include "defines.svh"
    `include "async_fifo_wr_seq_item.sv"
    `include "async_fifo_rd_seq_item.sv"
    `include "async_fifo_wr_sequence.sv"
    `include "async_fifo_rd_sequence.sv"
    `include "async_fifo_wr_sequencer.sv"
    `include "async_fifo_rd_sequencer.sv"
    `include "async_fifo_wr_driver.sv"
    `include "async_fifo_rd_driver.sv"
    `include "async_fifo_wr_monitor.sv"
    `include "async_fifo_rd_monitor.sv"
    `include "async_fifo_wr_agent.sv"
    `include "async_fifo_rd_agent.sv"
    `include "async_fifo_scoreboard_new.sv"
    `include "async_fifo_subscriber.sv"
    `include "async_fifo_virtual_sequencer.sv"
    `include "async_fifo_env.sv"
    `include "async_fifo_virtual_sequence.sv"
    `include "async_fifo_test.sv"
    
endpackage
